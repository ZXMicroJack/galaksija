XlxV38EB    fa00    2297(v׬ [�1CT =���2>hv+qS�|j������R� p�pC��oRe$���xm�b���בH�fr�"ʣ_�&�W��1nz��~W�F��7B���<Z�"�������K���16ϓM����{q�J��#�[��{Y	p����U�S��[�z���:�Ծxj/�k�� '�p�,��#;������l�Of��	=}��v+$I��)�C�[���8p��g�+(�K�r[���8����&�������L�,X��7��a8^���+*�6g�	Q�3_��m�9{(�:m��T!M���;~�QS�k��k ӢI~�k���%#������w��?h.��b#�M�n:7j
�iR[d?�s��PD��Y�^���Kâ�3��ξD�(�U%#r����(�&ÿ?�X�u���el��n�۔��k<���S�c�n�ٮ����׽R�]��d鼓5��𼟃���bs��D�<��Ы[�'�(W�sS"�]=M6-B5x�x͹	��j���E���b�"�2R��_�󀮬!  ���Y�ۍ�c���i��n�f_�8�$ ���t��Z*�}��}��V�!������e26A+���-�,Z
����(��M��Kk��%@�����'l�"H���bq��XW��C�]�ø#��jt���"��?�fq�_Syd�N��Y�bJg����F⶞@����H���	,v�d��'��-(+��ECʑe=�^���Q�'UۃKݑ��,0���h��|!��Z' cwmz4/�@��0>dRm���J���\tY�fv�'&���K��7��i�NѼ�,�'�3�0�-��3�qf��pޡq��x1>����[�>�2���н"����h�I+�t�x_��$=3�����aGyi(hМb!yM'c�(�@�Q�?�C����FQ�R`e�"U0她�~^C��p&O�O�ب��¹��O���C}�7͏0	ո ����<�������p�P�kc�ע�d��A�f���C�������1ͺc��#�U;�Z���A��Ü�����u��j���Q�_VJ��y\��M���5�� +�AA�����ڮ�Οa��b�EElj�"c1b�i8����{6qY�F,J��h[�i	���Z��6�D���Y�/.�����LIH>o^����3���	�l� @4�����q��޽@3<�H�a�f?Z7ؑ*�TKŲ��R��UD�`�~Jgi�S�&6F #���h�A�x���t����!| 5մ���m��x%Z��1B�L� + AMa������ q2��ˋ�55�pSx������}{Z�v>Y�:��cJ��h���Tb�2�e
�e��;���d���b�r���t���2,�M�'}�h(�� �=hX�7~�1� ء��[͓�$�K�&{{n ��Ļ�8��w�9/��I j��\=�dDM ;�4�)�9���	�<�̤꼗I#H�$��k]�Z����-f<:�K}8����f5�}���07B�Tq&:�z@����{��]\����^l��@��Ө�c6Uy7�64�7���A�w���K�Y���cj�<�oh�4������Q�M����r[(�?1ʫ&΁�c�nag��7��J_��>2�� 7;|�� �&ί{f�9:8u��b�a���V%��Dsg��ꮄi���:�Xv��U��"9�8�e�sѪҊE&K��D�A�u���Š=Z��?Q-�/���hL����8�m��5��،_���������͛��x�C� ���X�y�򡚯�4������˟5)��He�=�k�괰��]��֫x���R�5L��Mmc���d�7=�M��{������b�}N1-"�Y);�W*��O޹xC���e�Lu�85����{�'N�InGY���+��!+}g������/��W���
֝���X:z���^�^�j�0J�}Z<�&��0�<���_��,��%^>�A��Ĺ3�ל�8���
��P��� ڮwz�L{H�`�O҅}�u���Rh��\���rw��yE��'�S'D��82�_�z��9�����P��b�"2�N���ΠI�+��>M�v�U�t�]��P
���r.��܆%�����V�"6��H�*3����8�Kۢ��̈Xb���B����}��w�a���9�j>�� ^e��P��0����85{��~���*,�u[��3�e�����h��X�w�|�=s���*X��
ɐ�L��2��^�0:"}����xL�� ���Yr[�#<��Q�2!x�}��&9������1����½�R,��7��,E�iQ^�kl8�3�E�0�5��5�{�n������N'�e0��|��O�M��7��Y���N*�j�ٷr�]w��`� ����ו�kC0�6�#��	C��l.ζ?u��u�Hpx�����_ħ0Ȋ�7���>2�{2�5%���2O��H�[�/�#[%	��B��M��H�&�hfY�?�+���dU��_e�Mڞ����iw˄mںH`) m-.F�7�؎�r���H���>�p_p��Č����米��}��8����;��	S��)����i�����	�CDu�.�$��խ�"��3���ݼ?�ﳘ&��[ MW#�LJkH
V��czSG�?��u�C�yB �\UY�9˭�ܺU��\�(/!zDyGw�x��ߘI[�F}�MTq���Y�Ci�.Q�A�1��e���ΛyN�����\ �zS�y�j��;�n+�p^g�f���(сm��=CU̔������O�W�z�m��O�ko�A��H�����>��-��t�l��d���Y���2v��qYnfEX䏛�r�[
�c�	��5����-[�~
���3!����Yi�D��4�.c0�f�o�.�������5�=���H�.�
�}$2�`�u���a+�<��e��Ŝ_i�6`��,�٭nY�L�8f��G4q;̗��F�sJrT3�C�Jͣ��Ha
��8)�ea��~�kf3�>����6��0%7?T|X������׬�$0:QE@�P\�y��O]ԁ�5H�	\�㬑�EJ>ո@�"r{n]�l^H���,��HN%F.���9\�����ɔ[�F��bA>.���$�B�2�'Zwu�n�a^�l�<!����B�����t�t�V�M��E�^ ~�8�6��Fy{�`*�����ԏ�(�鼱�� �[��8���zF�m�)��}�!x1熷��a�n/���"��X�Y�U)x����!KH��D����k"�H	��_��{�e���g"N9.f$	��3K��@4zn�:-��YJ�>�9����0*�a��xE�Xy-/�g��[<w���n£�}O�)��WHr��:�b�y^��x�Gr.�Z�q[%<E�H,(�:=��Z�!C6�>P�y�O�ݎ=��������S�K�"�H�M�TPn
�Xv�>{�i#�����>���.s��$$�,�R�߆��HN4�Dze�T�I�"�l*8�ʄݯ�0O����;�O�,}���p
<������Gv��t2�f��.�te�Q
c�x�vMS�~�UJt�������}��׽�g�n�P�lv�!�y�D͠�����T�5���� ��d����.q޳��Z�|���U�Ƒ�=-g��=����"L�5� :�8!)�^'E�*���qV�eZ����ro+��=64�b��vR=H��R�{n�d�>�.�"X���7$ɷs�>���}���K ��>��G���.�S�6�{-��z��^�xY�7_�l����ݱ���^�ȹ���N��8M���vt�vVt4ї�.��XN����<�]���'�f��@�SJ������Cd��H���/�Bk �-�s/5b�Y����	�Bڢ��d,�ɘBDAfs&��Y�>P�#�?��%^r0=�-�?�yjFE��u�C{ڍ�%�7�#r���^�Eo4~�O�T&���<�.fG|Wm��edǇV�	� ư&a��&��
��)#���DEc��t��H�	x��͓kX�Ex����kj���!5_i�"}'%P'��7N�r�!]g��r�6:��'����Z"����݂B��Q���H�)r��sQ��Cǲl��K܇���<�n�ka�����&��n/��x)ёF�F�&�t�����Y�>����yD7�J��Q���+�6Y��@���Z���
C�E��j@��)�C��8��F>,J1J_���od���S(�_�矎)�p�[�n�i`�f�J��cյ��}�~ ����{
��GN}����Uż�b��#���&��I+�wZ �=�!2���=�w��v/q&���:j�,����༳�����Q��Ueb�נ�����Z���;a�f�%��{D�$)R����٩�ړ�T͂�S�ٹFz��=��� /���2��3}>�s�p��m2B��?/N��5�����ږX�}�ǔl�--r�7p4"E\�L��CV+5o��r3ݴ�d���ɦ�Vi������ㄆ���LM���}�;.�1{����_`���e�������h��P#y�C��D}��n:�YW|�.T/R�V�1����J�3Z�yj�e�e_$�
r�e@Z�q�7�K2��I��TP�%��8�����Q/�C{M�K\bZA��Q�J�	�5��Ϧ������W�S�;���L�aѺ��e�[ ����SP������R�r*�����]��B��Q���L��T�fA-���F�����Z܊�D��ep$.�%�ö�?;�@ӄ�Ќ&Rӿ[��y�"����f?��
��+4�8�a��}y�Wc�..�{����R�v�_ag{��������1SȦ«y4���ȁH�5
,���DD��U�&�����Z#r�t+���T�+��r�놽&�kS��uͨy#�S�u�t�`G���,�ή�PP)V"�ʰ5 �X�H�xr	q��a����ڎ(L�?*��D�&ð]: M�#��N���j��c�	na�v�����7���`����|�����/E^��]�d���e�#X���#$�Sv�x<�(�<����:�#�Pz��Q}U5,z��]�~���%�'�j���x��v�X'S�QSj4�{5I)?{��g)X�A���q�~Jo�ރ�)���uݗ�k�/�ѻE��v��[�\� �%�A������D�����C&��VA�pB�#�1i��cw���>�ȤZS;y�H_��B5�Q��idR��9V"O��Xv������h�)|3|[��2?2���}3��20�ɧ�����R��1��|�
:ϷC��N�Vv��/����Q���3u>RYe;��W�p8��f͡:L	�ʠs��7Ti����h�+�H
f�˝� �	;a�7h�tm��,ҍ4�W=�B�XbU�b�=w��W�����e��Fc�^~�*��%������Y��W.�	N����ǟ�.R�,&��&��h��T�8�֟�g.ōR6!\�r�3ɽZ����B.���	���a3$���l$���\4~����!�Z����>0�B���|�T)4�xG��&�ҵ�A�8nH�n^9�j�{?�νT��u�:����'u{�	,G_�Qk1���D�u��$0�6����w
"�E�6b���IngQ"��۽Ь�5+L&�[�^����}�T�&���#��[�J�6�Vd���D�M��rs��?�C��o�ӍO�Ӽ�����+�JVͩ��K�a�#�2'����0wH�*�׉�y7AX:�;��[4JA�&8и)��v�BEΞ`�jC-W�' v�=������?����=��B3 G��S�\�TY`�^�MJw@��W����z�j�w��\�!�)h���88��&& 2���C�8�6>�!"L��O��6ˉuP�Ϧ���!_�"��܊n�g+�B[\1 �֏=4�p��ޘ�����f#� C���Gh�VUc�M��4�𮁵��Qw�e̗�R���CH!��Q�y�����#!��\�'����q��*�upV�����B|��=Juw�d�G�#���x<zu�^#����Y���3�V���Z��bҒN����y-��ƨ�1�i}�=����-�\���JK�E�4@���4I��,�>A��^�Ĝ1`���+ú�LBd��a��~�����Pp^�1��]I�����1��^�.�J/K.\�V$T�m�ּ�`�!�}b��݃תH��,��!�p�M�q���yVZU0V�.��F�y��DK���a!�.-�P��R��N��D�;H��6�8P�_���\6�}�q�6�
ѳR+Y[?d��Uڧ͵Vwn{|K����
G481V60��W���.��_�����F�Ǝ�l�뛲]���Ak0��_�T�7�)�3�d�zS_�O�@ჱ�\��iU���*�l�A͙�B����C�U�{٩��>bGT�J� $�N��g3iu�K��e܎n��H�6w�	����B&e	"�%t��'�*E�����ۂt��"Ф��#z��L��͒Pk���!�Xͅ.����Cq�]��;r~�%J�u��S���.M~5��V��wsz/��.�Xt�#2ȿ�I��,{0z�Ae�/��*Qby��o4��Y��yO���q��W���KX����7��dX�K�'m�ފ��v�;4tn�d���-�vD�҂s���c`�W���	Y��H�Q l1�q�+z����Eaj%d/��-��������K��ﳏ$��n���O@>�kZ�_���Ṇ��E)��-G�&�t�`=�Z�ݫ�X��`��V�o�-P:��y�*n��<�^���\<`�S���q��餇D��r+o��8���L�1����a��X�ѣ�6�2��������Қ��_��B�	t�|���Y���x٭^<{kk��/B/���=�������M�b�����Y�*�a��%3U1;Pki2�����Ɇ�5�p�:>YN/�2_S�bB�d] �`D�T
K3p��y9�,-�����ˋHX�c�����9���m��/#K���������zU��?k�1-�_�
GQ�@���1���Bb���\�.�6_�oTT��ל�|����(]rϔ�ył��4���n%6C�.�]�W�(V��N�m>t��3��)m��/$�
����	�ܧX�浵�G*��˝�u탂/Q���p��G�0�2��aʤU�]�Y�f�X�j(��2D�0� ���(��\������}��}���	(�T�t��M�PQ���v�c�oK�p����W?!?H�	���/*��s���I�!�q�p_9A���f�h2C5�1��)�3�fUj����Ө/#,Z�>$5:UNz|`U%M$�cE7�Tͣ�h����Jg�c̔|;�n�_�x)]y�qJtr5�X��P�pf=/L)���$(L�V�sQ3ZF�:��r[%U�cD�=�</���|��-�b�~[I���i���o~�yJ�4��7�ֺ�/20�;w�F;	��?��.�!!/vBr���n�.U�㾄�"��95NH�|����x�;�����*M���.<�g\�����hm��5J��][~�s�G�	�K�U!��,(�ր��(zp%W��hD�E?�.Z!���.K�$�53W���T^9*k'ih����h����>c�J�sP�:2���S?�Ii�կ8�}Rh���Ҙ�%�Q@LRp��cסv�F�S�p}_)�,n_l<�AY1���Qr8�����Bt��o������,�SEY�{��M�B'8�z=}X|��`Vnۧ��%(؃j��}r7���(�Чm\/é��G��3��R����'�D���I�*���8;����U)�����Մ��%)/kOn�a�P��쇸���8����?`�n?�B�r���h�=N:$F�D]ceMP�@�G9]�Z�~�Y���	��s���)�ގ�-�D{����[�}!�����8Y�3'�� �����4��:�1E؅GR=[x��-vT$������덗	x��@� ��]�z�54^���B�:�zp@�]���+֯�|ff���ћ_O��[�jVn�^��3jn;��;�ĊrC3h�E��?���Gv�9n^&���m��~vQ�	oS"je��JE㇉$���@(۠3��>�
�8F�3�yiHNp�]�P 9xiH�c��^�Ρ!:v�B�*.���k��M��K2�W�#����|p����|[A�W�`%`�KS���3Ț�ë-��{Ͻ���d�JƳ����u�c'[���������*�d!���@Ūʢ�h8��������f�z*Y�����ʽ9��b�*ݿ	�@�qK;�K�� ��&�e�Ԉ�s6C��&]S	U�-�^S�^��W�El%�.��� hKq�2q�iN��cL�6<�\�j��z��R��_Y�o���ºS��������t��/����~x&[�Iz�yƬ��(xS�NXj�0|ٶ`A�b�p���>��_���#�u����!����]�ͬ&sg;�旡pТm���
�wd<��G���2T�q_�yƅ�o���E��$����2�D�y����C�3u1ߨG�v_�<�`Ό��K_=�?�NT�XlxV38EB     761     14c�c0^A�U�Ni�x��
�{���Uy��%G*8W۸�E)�����my�ۨ���*r���]5E|�~��+j���Abe]��]���<�=��*�R�.J��hY�R��z}��cÚ??��|��Z!dQ�qQHJ2&F�]�Kd>�^Y����cF�[�,��HyS��b]l�I�Xlm������rxW�{8apzb�Ӆ'���T����H�y��:�va�<��$gŵˉk+!������-]�۲��>�-��SL�\�8bC>�г/ �)��fto��e6U5^��R�v�~ �bV�"��HoGW{й[(�$�ˣa���